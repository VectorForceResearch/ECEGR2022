--------------------------------------------------------------------------------
--
-- LAB #5 - Memory and Register Bank
--
--------------------------------------------------------------------------------
LIBRARY ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity RAM is
    Port(Reset:	  in std_logic;
         Clock:	  in std_logic;
         OE:      in std_logic;
         WE:      in std_logic;
         Address: in std_logic_vector(29 downto 0);
         DataIn:  in std_logic_vector(31 downto 0);
         DataOut: out std_logic_vector(31 downto 0));
end entity RAM;

architecture staticRAM of RAM is

   type ram_type is array (0 to 127) of std_logic_vector(31 downto 0);
   signal i_ram : ram_type;

begin

  RamProc: process(Clock, Reset, OE, WE, Address) is

  begin
    if Reset = '1' then
      for i in 0 to 127 loop
          i_ram(i) <= X"00000000";
      end loop;
    end if;

    if falling_edge(Clock) then
  -- Add code to write data to RAM
  -- Use to_integer(unsigned(Address)) to index the i_ram array
      if WE = '1' then
          for i in 0 to 127 loop
              i_ram(i) <= DataIn(i);
              -- found doc that this might work: RamProc(address) := DataIn(i);
          end loop;
      end if;

      if OE = '0' then
          for i in 0 to 127 loop
              DataOut(i) <= i_ram(i);
              -- found doc that this might work: DataOut(i) <= RamProc(Address);
          end loop;
      end if;
    end if;

  -- Rest of the RAM implementation

  end process RamProc;

end staticRAM;


--------------------------------------------------------------------------------
LIBRARY ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity Registers is
    Port(ReadReg1: in std_logic_vector(4 downto 0);
         ReadReg2: in std_logic_vector(4 downto 0);
         WriteReg: in std_logic_vector(4 downto 0);
         WriteData: in std_logic_vector(31 downto 0);
         WriteCmd: in std_logic;
         ReadData1: out std_logic_vector(31 downto 0);
         ReadData2: out std_logic_vector(31 downto 0));
end entity Registers;

architecture remember of Registers is
  component register32
  	    port(datain: in std_logic_vector(31 downto 0);
             enout32,enout16,enout8: in std_logic;
             writein32, writein16, writein8: in std_logic;
             dataout: out std_logic_vector(31 downto 0));
  end component;

begin
    -- Add your code here for the Register Bank implementation

    RegProc: process(WriteCmd) is

    end RegProc;

end remember;

----------------------------------------------------------------------------------------------------------------------------------------------------------------
